version https://git-lfs.github.com/spec/v1
oid sha256:58361591fdea63cbecebff577e43e51a41426b7e7f758cd733faf844bdd16bc3
size 18658
