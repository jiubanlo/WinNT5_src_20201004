version https://git-lfs.github.com/spec/v1
oid sha256:8405adb317f48613fb49d5900081954ce72cfcfba36cd7338ce4b77053a547ff
size 19351
