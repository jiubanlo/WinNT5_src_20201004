version https://git-lfs.github.com/spec/v1
oid sha256:f5ca3ac3a250837e27f6228a1c00b519e8f0c7a6e5e31ddc5a6077489cba19ea
size 76542
